module ShiftDecoder2(input Shift_Left, input Shift_Right, input BFE, input [3:0] SL, input [3:0] SR, output [3:0] X, output [3:0] Y, output [3:0] Z);

assign X[3] = (Shift_Left|BFE)&SL[3];
assign X[2] = (Shift_Left|BFE)&SL[2];
assign X[1] = (Shift_Left|BFE)&SL[1];
assign X[0] = (Shift_Left|BFE)&SL[0];

wire [3:0] sum;

assign sum = SL+SR;

assign Y[3] = (Shift_Right&SR[3])|(BFE&sum[3]);
assign Y[2] = (Shift_Right&SR[2])|(BFE&sum[2]);
assign Y[1] = (Shift_Right&SR[1])|(BFE&sum[1]);
assign Y[0] = (Shift_Right&SR[0])|(BFE&sum[0]);

assign Z[3] = BFE&SR[3];
assign Z[2] = BFE&SR[2];
assign Z[1] = BFE&SR[1];
assign Z[0] = BFE&SR[0];



endmodule