module Decoder ()

input [4..0] ir;



assign stp = !ir[4] & !ir[3] & !ir[2] & !ir[1] & !ir[0];
assign adr = !ir[4] & !ir[3] & !ir[2] & !ir[1] &  ir[0];
assign adm = !ir[4] & !ir[3] & !ir[2] &  ir[1] & !ir[0];
assign adi = !ir[4] & !ir[3] & !ir[2] &  ir[1] &  ir[0];
assign sbr = !ir[4] & !ir[3] &  ir[2] & !ir[1] & !ir[0];
assign sbm = !ir[4] & !ir[3] &  ir[2] & !ir[1] &  ir[0];
assign sbi = !ir[4] & !ir[3] &  ir[2] &  ir[1] & !ir[0];
assign mlr = !ir[4] & !ir[3] &  ir[2] &  ir[1] &  ir[0];
assign mlm = !ir[4] &  ir[3] & !ir[2] & !ir[1] & !ir[0];
assign xsl = !ir[4] &  ir[3] & !ir[2] & !ir[1] &  ir[0];
assign xsr = !ir[4] &  ir[3] & !ir[2] &  ir[1] & !ir[0];
assign bbo = !ir[4] &  ir[3] & !ir[2] &  ir[1] &  ir[0];
assign bfe = !ir[4] &  ir[3] &  ir[2] & !ir[1];
assign jmr = !ir[4] &  ir[3] &  ir[2] &  ir[1] &  ir[0];
assign jmp = !ir[4] &  ir[3] &  ir[2] &  ir[1] &
assign ldi =  ir[4] & !ir[3] & !ir[2];
assign sta =  ir[4] & !ir[3] &  ir[2];
assign ldr =  ir[4] &  ir[3] & !ir[2] & !ir[1] & !ir[0];
assign sti =  ir[4] &  ir[3] & !ir[2] & !ir[1] &  ir[0];
assign psh =  ir[4] &  ir[3] & !ir[2] &  ir[1] & !ir[0];
assign pop =  ir[4] &  ir[3] & !ir[2] &  ir[1] &  ir[0];