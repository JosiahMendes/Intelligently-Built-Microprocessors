module halfAdderNoC(input A, input B, output S);

assign S = A ^ B;

endmodule