
module OR15(input A,B,C,D,E,F,G,H,I,J,K,L,M,N,O, output Cout);

assign Cout = A|B|C|D|E|F|G|H|I|J|K|L|M|N|O; 

endmodule